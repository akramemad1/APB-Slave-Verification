package APB_Coverage_Class_pkg;


class APB_Coverage_Class;





endclass //APB_Coverage_Class

    
endpackage